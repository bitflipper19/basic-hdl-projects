// 4-bit carry look ahead adder [Generate and Propagate focussed]

module cla4bit (
    output [3:0] SUM,
    output carry,
    input [3:0] A, B,
    input C0
);
    
endmodule