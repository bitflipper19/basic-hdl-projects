module ic_7483(

);